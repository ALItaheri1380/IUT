module top;
	reg [15:0] a;
	reg [2:0] b;
	wire [4:0] out;
	log g1(a , b , out);
	
	initial
	begin
		#100{a , b} = 19'b0000000000011100011;//28 ->3
		#100{a , b} = 19'b0000000000001110100;//14 ->4
		#100{a , b} = 19'b0000000000111110010;//62 ->2
		#100{a , b} = 19'b0000000000000011010;//3 ->2
		#100{a , b} = 19'b0000000000001000011;
		#100;
	end
endmodule
