module not_gate(a , o);
   
   input a;
   output o;
   nor(o , a , a);

endmodule
